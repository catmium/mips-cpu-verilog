module pc ();



endmodule