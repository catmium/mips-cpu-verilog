module alu ();

endmodule